module IF_ID_Register(reset,
                      clk,
                      i_pc_4,
                      i_instruction,
                      i_flush,
                      o_pc_4,
                      o_instruction);
    input reset;
    input clk;
    input i_flush;
    input [31:0] i_pc_4;
    input [31:0] i_instruction;
    
    output reg [31:0] o_pc_4;
    output reg [31:0] o_instruction;
    
    always @(posedge reset or posedge clk) begin
        if(reset) begin
            o_pc_4 <= 32'b0;
            o_instruction <= 32'b0;
        end
        else begin
            if(i_flush) begin // a 'nop' command is generated by hazard unit
                o_instruction <= 32'b0;
            end
            else begin
                o_instruction <= i_instruction;
            end
            o_pc_4 <= i_pc_4;
        end

    end
endmodule
