module ID_Forward(
    
);

endmodule