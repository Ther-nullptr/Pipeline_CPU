`timescale 1ns / 1ps
module InstructionMemory(i_address,
                         o_instruction);
    
    input [8:0] i_address;
    output reg [31:0] o_instruction;
    always @(*)
        case (i_address)
            9'd0:    o_instruction   <= 32'h20100000;
            9'd1:    o_instruction   <= 32'h20050000;
            9'd2:    o_instruction   <= 32'h20060001;
            9'd3:    o_instruction   <= 32'h8ca80000;
            9'd4:    o_instruction   <= 32'h2009000a;
            9'd5:    o_instruction   <= 32'h11090003;
            9'd6:    o_instruction   <= 32'h20a50004;
            9'd7:    o_instruction   <= 32'h22100001;
            9'd8:    o_instruction   <= 32'h08000003;
            9'd9:    o_instruction   <= 32'h20a50004;
            9'd10:    o_instruction  <= 32'h20b20000;
            9'd11:    o_instruction  <= 32'h20060001;
            9'd12:    o_instruction  <= 32'h20110000;
            9'd13:    o_instruction  <= 32'h8ca80000;
            9'd14:    o_instruction  <= 32'h2009000a;
            9'd15:    o_instruction  <= 32'h11090003;
            9'd16:    o_instruction  <= 32'h20a50004;
            9'd17:    o_instruction  <= 32'h22310001;
            9'd18:    o_instruction  <= 32'h0800000d;
            9'd19:    o_instruction  <= 32'h22040000;
            9'd20:    o_instruction  <= 32'h20050000;
            9'd21:    o_instruction  <= 32'h22260000;
            9'd22:    o_instruction  <= 32'h00123820;
            9'd23:    o_instruction  <= 32'h0c000042;
            9'd24:    o_instruction  <= 32'h20500000;
            9'd25:    o_instruction  <= 32'h00108f00;
            9'd26:    o_instruction  <= 32'h00118f02;
            9'd27:    o_instruction  <= 32'h00109600;
            9'd28:    o_instruction  <= 32'h00129702;
            9'd29:    o_instruction  <= 32'h00109d00;
            9'd30:    o_instruction  <= 32'h00139f02;
            9'd31:    o_instruction  <= 32'h0010a400;
            9'd32:    o_instruction  <= 32'h0014a702;
            9'd33:    o_instruction  <= 32'h3c164000;
            9'd34:    o_instruction  <= 32'h22d60014;
            9'd35:    o_instruction  <= 32'h200d2710;
            9'd36:    o_instruction  <= 32'h200e4e20;
            9'd37:    o_instruction  <= 32'h200f7530;
            9'd38:    o_instruction  <= 32'h200c0100;
            9'd39:    o_instruction  <= 32'h22240000;
            9'd40:    o_instruction  <= 32'h0c0000a2;
            9'd41:    o_instruction  <= 32'h8ed70000;
            9'd42:    o_instruction  <= 32'h02ed5822;
            9'd43:    o_instruction  <= 32'h1d600001;
            9'd44:    o_instruction  <= 32'h08000026;
            9'd45:    o_instruction  <= 32'h200c0200;
            9'd46:    o_instruction  <= 32'h22440000;
            9'd47:    o_instruction  <= 32'h0c0000a2;
            9'd48:    o_instruction  <= 32'h8ed70000;
            9'd49:    o_instruction  <= 32'h02ee5822;
            9'd50:    o_instruction  <= 32'h1d600001;
            9'd51:    o_instruction  <= 32'h0800002d;
            9'd52:    o_instruction  <= 32'h200c0400;
            9'd53:    o_instruction  <= 32'h22640000;
            9'd54:    o_instruction  <= 32'h0c0000a2;
            9'd55:    o_instruction  <= 32'h8ed70000;
            9'd56:    o_instruction  <= 32'h02ef5822;
            9'd57:    o_instruction  <= 32'h1d600001;
            9'd58:    o_instruction  <= 32'h08000034;
            9'd59:    o_instruction  <= 32'h200c0800;
            9'd60:    o_instruction  <= 32'h22840000;
            9'd61:    o_instruction  <= 32'h0c0000a2;
            9'd62:    o_instruction  <= 32'h8ed70000;
            9'd63:    o_instruction  <= 32'h02ed5822;
            9'd64:    o_instruction  <= 32'h0560ffe5;
            9'd65:    o_instruction  <= 32'h0800003b;
            9'd66:    o_instruction  <= 32'h23bdfffc;
            9'd67:    o_instruction  <= 32'hafbf0000;
            9'd68:    o_instruction  <= 32'h20940000;
            9'd69:    o_instruction  <= 32'h20d50000;
            9'd70:    o_instruction  <= 32'h20b60000;
            9'd71:    o_instruction  <= 32'h20f70000;
            9'd72:    o_instruction  <= 32'h20100300;
            9'd73:    o_instruction  <= 32'h22040000;
            9'd74:    o_instruction  <= 32'h20c50000;
            9'd75:    o_instruction  <= 32'h20e60000;
            9'd76:    o_instruction  <= 32'h0c000071;
            9'd77:    o_instruction  <= 32'h20100000;
            9'd78:    o_instruction  <= 32'h20110000;
            9'd79:    o_instruction  <= 32'h20120000;
            9'd80:    o_instruction  <= 32'h1214001c;
            9'd81:    o_instruction  <= 32'h00104080;
            9'd82:    o_instruction  <= 32'h00114880;
            9'd83:    o_instruction  <= 32'h02e96020;
            9'd84:    o_instruction  <= 32'h02c86820;
            9'd85:    o_instruction  <= 32'h8d8e0000;
            9'd86:    o_instruction  <= 32'h8daf0000;
            9'd87:    o_instruction  <= 32'h15cf000c;
            9'd88:    o_instruction  <= 32'h22abffff;
            9'd89:    o_instruction  <= 32'h162b0007;
            9'd90:    o_instruction  <= 32'h22520001;
            9'd91:    o_instruction  <= 32'h22b8ffff;
            9'd92:    o_instruction  <= 32'h0018c080;
            9'd93:    o_instruction  <= 32'h0313c020;
            9'd94:    o_instruction  <= 32'h8f110000;
            9'd95:    o_instruction  <= 32'h22100001;
            9'd96:    o_instruction  <= 32'h0800006c;
            9'd97:    o_instruction  <= 32'h22310001;
            9'd98:    o_instruction  <= 32'h22100001;
            9'd99:    o_instruction  <= 32'h0800006c;
            9'd100:    o_instruction <= 32'h0011c82a;
            9'd101:    o_instruction <= 32'h13200005;
            9'd102:    o_instruction <= 32'h2238ffff;
            9'd103:    o_instruction <= 32'h0018c080;
            9'd104:    o_instruction <= 32'h0313c020;
            9'd105:    o_instruction <= 32'h8f110000;
            9'd106:    o_instruction <= 32'h0800006c;
            9'd107:    o_instruction <= 32'h22100001;
            9'd108:    o_instruction <= 32'h08000050;
            9'd109:    o_instruction <= 32'h22420000;
            9'd110:    o_instruction <= 32'h8fbf0000;
            9'd111:    o_instruction <= 32'h23bd0004;
            9'd112:    o_instruction <= 32'h03e00008;
            9'd113:    o_instruction <= 32'h23bdfff4;
            9'd114:    o_instruction <= 32'hafb00008;
            9'd115:    o_instruction <= 32'hafb10004;
            9'd116:    o_instruction <= 32'hafb20000;
            9'd117:    o_instruction <= 32'h20110001;
            9'd118:    o_instruction <= 32'h20120000;
            9'd119:    o_instruction <= 32'h20010000;
            9'd120:    o_instruction <= 32'h1025001d;
            9'd121:    o_instruction <= 32'h20d00000;
            9'd122:    o_instruction <= 32'h20930000;
            9'd123:    o_instruction <= 32'hae600000;
            9'd124:    o_instruction <= 32'h1225001f;
            9'd125:    o_instruction <= 32'h00115080;
            9'd126:    o_instruction <= 32'h00124080;
            9'd127:    o_instruction <= 32'h020a6020;
            9'd128:    o_instruction <= 32'h02086820;
            9'd129:    o_instruction <= 32'h8d8c0000;
            9'd130:    o_instruction <= 32'h8dad0000;
            9'd131:    o_instruction <= 32'h158d0006;
            9'd132:    o_instruction <= 32'h22480001;
            9'd133:    o_instruction <= 32'h026a7820;
            9'd134:    o_instruction <= 32'hade80000;
            9'd135:    o_instruction <= 32'h22520001;
            9'd136:    o_instruction <= 32'h22310001;
            9'd137:    o_instruction <= 32'h08000095;
            9'd138:    o_instruction <= 32'h0012702a;
            9'd139:    o_instruction <= 32'h11c00005;
            9'd140:    o_instruction <= 32'h224fffff;
            9'd141:    o_instruction <= 32'h000f5080;
            9'd142:    o_instruction <= 32'h026a7820;
            9'd143:    o_instruction <= 32'h8df20000;
            9'd144:    o_instruction <= 32'h08000095;
            9'd145:    o_instruction <= 32'h00115080;
            9'd146:    o_instruction <= 32'h026a7820;
            9'd147:    o_instruction <= 32'hade00000;
            9'd148:    o_instruction <= 32'h22310001;
            9'd149:    o_instruction <= 32'h0800007c;
            9'd150:    o_instruction <= 32'h20020001;
            9'd151:    o_instruction <= 32'h8fb00008;
            9'd152:    o_instruction <= 32'h8fb10004;
            9'd153:    o_instruction <= 32'h8fb20000;
            9'd154:    o_instruction <= 32'h23bd000c;
            9'd155:    o_instruction <= 32'h03e00008;
            9'd156:    o_instruction <= 32'h20020000;
            9'd157:    o_instruction <= 32'h8fb00008;
            9'd158:    o_instruction <= 32'h8fb10004;
            9'd159:    o_instruction <= 32'h8fb20000;
            9'd160:    o_instruction <= 32'h23bd000c;
            9'd161:    o_instruction <= 32'h03e00008;
            9'd162:    o_instruction <= 32'h20080000;
            9'd163:    o_instruction <= 32'h1088001e;
            9'd164:    o_instruction <= 32'h20080001;
            9'd165:    o_instruction <= 32'h1088001e;
            9'd166:    o_instruction <= 32'h20080002;
            9'd167:    o_instruction <= 32'h1088001e;
            9'd168:    o_instruction <= 32'h20080003;
            9'd169:    o_instruction <= 32'h1088001e;
            9'd170:    o_instruction <= 32'h20080004;
            9'd171:    o_instruction <= 32'h1088001e;
            9'd172:    o_instruction <= 32'h20080005;
            9'd173:    o_instruction <= 32'h1088001e;
            9'd174:    o_instruction <= 32'h20080006;
            9'd175:    o_instruction <= 32'h1088001e;
            9'd176:    o_instruction <= 32'h20080007;
            9'd177:    o_instruction <= 32'h1088001e;
            9'd178:    o_instruction <= 32'h20080008;
            9'd179:    o_instruction <= 32'h1088001e;
            9'd180:    o_instruction <= 32'h20080009;
            9'd181:    o_instruction <= 32'h1088001e;
            9'd182:    o_instruction <= 32'h2008000a;
            9'd183:    o_instruction <= 32'h1088001e;
            9'd184:    o_instruction <= 32'h2008000b;
            9'd185:    o_instruction <= 32'h1088001e;
            9'd186:    o_instruction <= 32'h2008000c;
            9'd187:    o_instruction <= 32'h1088001e;
            9'd188:    o_instruction <= 32'h2008000d;
            9'd189:    o_instruction <= 32'h1088001e;
            9'd190:    o_instruction <= 32'h2008000e;
            9'd191:    o_instruction <= 32'h1088001e;
            9'd192:    o_instruction <= 32'h2008000f;
            9'd193:    o_instruction <= 32'h1088001e;
            9'd194:    o_instruction <= 32'h2009003f;
            9'd195:    o_instruction <= 32'h080000e2;
            9'd196:    o_instruction <= 32'h20090006;
            9'd197:    o_instruction <= 32'h080000e2;
            9'd198:    o_instruction <= 32'h2009005b;
            9'd199:    o_instruction <= 32'h080000e2;
            9'd200:    o_instruction <= 32'h2009004f;
            9'd201:    o_instruction <= 32'h080000e2;
            9'd202:    o_instruction <= 32'h20090066;
            9'd203:    o_instruction <= 32'h080000e2;
            9'd204:    o_instruction <= 32'h2009006d;
            9'd205:    o_instruction <= 32'h080000e2;
            9'd206:    o_instruction <= 32'h2009007d;
            9'd207:    o_instruction <= 32'h080000e2;
            9'd208:    o_instruction <= 32'h20090007;
            9'd209:    o_instruction <= 32'h080000e2;
            9'd210:    o_instruction <= 32'h2009007f;
            9'd211:    o_instruction <= 32'h080000e2;
            9'd212:    o_instruction <= 32'h2009006f;
            9'd213:    o_instruction <= 32'h080000e2;
            9'd214:    o_instruction <= 32'h20090077;
            9'd215:    o_instruction <= 32'h080000e2;
            9'd216:    o_instruction <= 32'h2009007c;
            9'd217:    o_instruction <= 32'h080000e2;
            9'd218:    o_instruction <= 32'h20090039;
            9'd219:    o_instruction <= 32'h080000e2;
            9'd220:    o_instruction <= 32'h2009005e;
            9'd221:    o_instruction <= 32'h080000e2;
            9'd222:    o_instruction <= 32'h20090079;
            9'd223:    o_instruction <= 32'h080000e2;
            9'd224:    o_instruction <= 32'h20090071;
            9'd225:    o_instruction <= 32'h080000e2;
            9'd226:    o_instruction <= 32'h3c154000;
            9'd227:    o_instruction <= 32'h22b50010;
            9'd228:    o_instruction <= 32'h012c4820;
            9'd229:    o_instruction <= 32'haea90000;
            9'd230:    o_instruction <= 32'h03e00008;
            default: o_instruction   <= 32'h00000000;
        endcase
endmodule
