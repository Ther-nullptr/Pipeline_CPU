`timescale 1ns / 1ps

module InstructionMemory(
    i_address,
    o_instruction
);

    input [31:0] i_address;
    output [31:0] o_instruction;

endmodule